/*	AND_2	*/
module	AND_2	( IN1, IN2, OUT );
input	IN1, IN2;			// Set input variable name 
output	OUT;				// Set output variable name
	and	U1	( OUT, IN1, IN2 );
endmodule
